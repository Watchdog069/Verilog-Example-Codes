//design code
module andgate(y,a,b);
	output y;
	input a;
	input b;
	assign y=a|b;
endmodule